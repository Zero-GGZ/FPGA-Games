/*=======================================================
Author				:				QiiNn
Email Address		:				ctlvie@gmail.com
Filename			:				showtank_app.v
Date				:				2018-05-12
Description			:				

Modification History:
Date		By			Version		Description
----------------------------------------------------------
========================================================*/

`timescale 1ns/1ns

module showtank_app
(	
	input 			clk,
	input 			clk_4Hz,
	input 			enable,
	input	[4:0]	start_x,
	input	[4:0]	start_y,
	input	[1:0]	start_dir,
	input			bul_state_feedback,
	output	reg 	[4:0]	x_rel_pos_out,
	output	reg 	[4:0]	y_rel_pos_out,		
	output	reg	[1:0]		tank_dir_out,
	output  reg				bul_sht
);

reg 	tank_state_reg;
reg		[3:0]	cnt;
//---------------------------------------------------
//initial coordinate generation

reg sample;
initial sample <= 1'b0;
//---------------------------------------------------
//moving
always@(posedge clk_4Hz)
begin
if(enable)
begin
	if(!sample)
		begin
		x_rel_pos_out <= start_x;
		y_rel_pos_out <= start_y;
		sample <= 1'b1;
		end
	//move upward and direction = 00
	if(start_dir == 2'b00)
	begin
		y_rel_pos_out <= y_rel_pos_out - 1'b1;
		tank_dir_out <= 2'b00;
		if (y_rel_pos_out == 0)
			y_rel_pos_out <= 12; 
	end

	//move downward and direction = 01
	if(start_dir == 2'b01)
	begin
		y_rel_pos_out <= y_rel_pos_out + 1'b1;
		tank_dir_out <= 2'b01;
		if (y_rel_pos_out == 12)
			y_rel_pos_out <= 0; 
	end

	//move left and direction = 10
	if(start_dir == 2'b10)
	begin
		x_rel_pos_out <= x_rel_pos_out - 1'b1;
		tank_dir_out <= 2'b10;
		if (x_rel_pos_out == 0)
			x_rel_pos_out <= 24; 
	end

	//move right and direction = 11
	if(start_dir == 2'b11)
	begin
		x_rel_pos_out <= x_rel_pos_out + 1'b1;
		tank_dir_out <= 2'b11;
		if (x_rel_pos_out == 24)
			x_rel_pos_out <= 0; 
	end
end
end

//---------------------------------------------------
//Shoot

always@(posedge clk_4Hz)
	cnt <= cnt + 1;
/*
always@(posedge clk)
begin
if(enable)
begin
	if (bul_state_feedback == 1'b0)
	begin
		if (cnt == 0)
			bul_sht <= 1'b1;
		else
			bul_sht <= 1'b0;	
	end
	else
	begin
		bul_sht <= 1'b1;
	end
end
end
*/

reg [10:0]	cnt;
initial cnt <= 0;
/*
always@(posedge clk)
begin
if(enable)
begin
	if (bul_state_feedback == 1'b0)
	begin
		bul_sht <= 0;
		cnt <= cnt + 1;
		if (cnt >= 20000)
		begin
			bul_sht <= 1;
			cnt <= 0;
		end
	end
	else
		bul_sht <= 1;
end
end
*/

always@(posedge clk)
begin
if(enable)
	begin
	bul_sht <= 1;
	end
else
	bul_sht <= 0;
end
endmodule